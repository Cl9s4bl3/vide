module lib

pub fn cd(args []string) int {
	println("Hello world!")
	return 0
}